* AD8056 SPICE model
* Description: Amplifier
* Generic Desc: Dual 300 MHz voltage feedback op amp
* Developed by: SMR/ADI
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (08/1997)
* Copyright 1997, 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*     distortion is not characterized
*
* Parameters modeled include:
*     closed loop gain and phase vs bandwidth
*     output current and voltage limiting
*     offset voltage (is static, will not vary with vcm)
*     ibias (again, is static, will not vary with vcm)
*     slew rate and step response performance
*     (slew rate is based on 10-90% of step response)
*     current on output will be reflected to the supplies
*     vnoise, referred to the input
*     inoise, referred to the input
*
* END Notes
*
* Node assignments
* 		 non-inverting input
*                | inverting input
*                | | positive supply
*                | | |  negative supply
*                | | |  | output
*                | | |  |  |
.SUBCKT AD8056   1 2 99 50 17

* input stage
*
q1 4 15 13 qn1
q2 5 2 14 qn1
i1 3 50 0.1
i2 50 99 0.1
r3 99 4 14.96
r4 99 5 14.96
r5 13 3 14.44
r6 14 3 14.44
cpole 4 5 26.61pf
cin1 1 98 2pf
cin2 2 98 2pf

* error stage

eos 1 15 poly(2) 30 98 92 0 3e-3 1 25e-9
gnoise1 98 1 33 98 1e-4
gnoise2 98 2 33 98 1e-4

* gain/bw stage

g1 99 9 poly(1) 5 4 0 0.067 0 0.022
g2 50 9 poly(1) 5 4 0 0.067 0 0.022
rgain1 99 9 53078
rgain2 50 9 53078
cgain1 99 9 71.42pf
cgain2 50 9 71.42pf
vlim1 99 18 2.46
vlim2 19 50 2.46
dlim1 9 18 d1
dlim2 19 9 d1

* vnoise stage
*

rnoise1 39 98 0.46e-3
vnoise1 39 98 0
vnoise2 31 98 0.56
dnoise1 31 39 dn
fnoise1 30 98 vnoise1 1
rnoise2 30 98 1

* inoise stage
*

rnoise3 32 98 0.166e-3
vnoise3 32 98 0
vnoise4 34 98 0.545
dnoise2 34 32 dn
fnoise2 33 98 vnoise3 1
rnoise4 33 98 1

* buffer stage

gbuf 98 12 9 98 1e-2
rbuf 98 12 100

* reference stage

eref1 98 0 poly(2) 99 0 50 0 0 0.5 0.5
eref2 97 0 poly(2) 1 0 2 0 0 0.5 0.5

* common mode rejection
*

ecm1 96 0 98 97 23809
rcm2 96 95 23809
rcm1 95 94 1
lcm1 94 0 3.79e-6
ecm2 93 0 95 0 3332
rcm3 93 92 3332
rcm4 92 89 1
lcm2 89 0 0.53e-6

* output current reflected to supplies
*

fcurr 98 40 vout 1
vcur1 26 98 0
vcur2 98 27 0
dcur1 40 26 d1
dcur2 27 40 d1

* output stage

vo1 99 90 0
vo2 91 50 0
fout1 0 99 poly(2) vo1 vcur1 -5.4e-3 1 -1
fout2 50 0 poly(2) vo2 vcur2 -5.4e-3 1 -1
gout1 90 16 12 99 1
gout2 91 16 12 50 1
rout1 16 90 1
rout2 16 91 1
vout 16 17 0
viclmp1 12 20 0.703
viclmp2 21 12 0.703
diclmp1 16 20 d1
diclmp2 21 16 d1
.model qn1 npn(bf=1e5)
.model d1  d()
.model dn  d(af=1 kf=1e-8)
.ends ad8056






